-------------------------------------------

-- Construa um circuito que lê NUM_SWITCHES chaves como um número binário e NUM_BUTTONS como uma exponenciação de base	
-- binária (e.g. 2 botões apertados -> 2**2 = 4) e multiplica esses dois valores, mostrando o resultado nos SSDs.	
-- Esse exercício deve ser completamente genérico.

-------------------------------------------

library ieee;

use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.math_real.all;
use work.own_Library.all;

-------------------------------------------

entity Laboratorio_06_02 is
	generic (
	
	);
	
	port (
	
	);
end entity;

-------------------------------------------

architecture Laboratorio_06_02 of Laboratorio_06_02 is
	
	begin
		
end architecture;

